//
// Copyright (C) 2024, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
//

module tst_dout_xclk
(
	//--------------------------------
	// register clock domain
	//--------------------------------
	input   clk_reg,
	input   rst_reg,
	input   test_en_reg,
	output  [47:0] r00_smp_reg,
	output  [47:0] r00_err_reg,
	output  [47:0] r00_idl_reg,
	output  [15:0] r00_lat_reg,
	output  [47:0] r01_smp_reg,
	output  [47:0] r01_err_reg,
	output  [47:0] r01_idl_reg,
	output  [15:0] r01_lat_reg,	
	output  [47:0] r02_smp_reg,
	output  [47:0] r02_err_reg,
	output  [47:0] r02_idl_reg,
	output  [15:0] r02_lat_reg,
	output  [47:0] r03_smp_reg,
	output  [47:0] r03_err_reg,
	output  [47:0] r03_idl_reg,
	output  [15:0] r03_lat_reg,
	output  [47:0] r04_smp_reg,
	output  [47:0] r04_err_reg,
	output  [47:0] r04_idl_reg,
	output  [15:0] r04_lat_reg,
	output  [47:0] r05_smp_reg,
	output  [47:0] r05_err_reg,
	output  [47:0] r05_idl_reg,
	output  [15:0] r05_lat_reg,	
	output  [47:0] r06_smp_reg,
	output  [47:0] r06_err_reg,
	output  [47:0] r06_idl_reg,
	output  [15:0] r06_lat_reg,
	output  [47:0] r07_smp_reg,
	output  [47:0] r07_err_reg,
	output  [47:0] r07_idl_reg,
	output  [15:0] r07_lat_reg,
	output  [47:0] r10_smp_reg,
	output  [47:0] r10_err_reg,
	output  [47:0] r10_idl_reg,
	output  [15:0] r10_lat_reg,
	output  [47:0] r11_smp_reg,
	output  [47:0] r11_err_reg,
	output  [47:0] r11_idl_reg,
	output  [15:0] r11_lat_reg,	
	output  [47:0] r12_smp_reg,
	output  [47:0] r12_err_reg,
	output  [47:0] r12_idl_reg,
	output  [15:0] r12_lat_reg,
	output  [47:0] r13_smp_reg,
	output  [47:0] r13_err_reg,
	output  [47:0] r13_idl_reg,
	output  [15:0] r13_lat_reg,
	output  [47:0] r14_smp_reg,
	output  [47:0] r14_err_reg,
	output  [47:0] r14_idl_reg,
	output  [15:0] r14_lat_reg,
	output  [47:0] r15_smp_reg,
	output  [47:0] r15_err_reg,
	output  [47:0] r15_idl_reg,
	output  [15:0] r15_lat_reg,	
	output  [47:0] r16_smp_reg,
	output  [47:0] r16_err_reg,
	output  [47:0] r16_idl_reg,
	output  [15:0] r16_lat_reg,
	output  [47:0] r17_smp_reg,
	output  [47:0] r17_err_reg,
	output  [47:0] r17_idl_reg,
	output  [15:0] r17_lat_reg,	
	output  [47:0] r20_smp_reg,
	output  [47:0] r20_err_reg,
	output  [47:0] r20_idl_reg,
	output  [15:0] r20_lat_reg,
	output  [47:0] r21_smp_reg,
	output  [47:0] r21_err_reg,
	output  [47:0] r21_idl_reg,
	output  [15:0] r21_lat_reg,	
	output  [47:0] r22_smp_reg,
	output  [47:0] r22_err_reg,
	output  [47:0] r22_idl_reg,
	output  [15:0] r22_lat_reg,
	output  [47:0] r23_smp_reg,
	output  [47:0] r23_err_reg,
	output  [47:0] r23_idl_reg,
	output  [15:0] r23_lat_reg,
	output  [47:0] r24_smp_reg,
	output  [47:0] r24_err_reg,
	output  [47:0] r24_idl_reg,
	output  [15:0] r24_lat_reg,
	output  [47:0] r25_smp_reg,
	output  [47:0] r25_err_reg,
	output  [47:0] r25_idl_reg,
	output  [15:0] r25_lat_reg,	
	output  [47:0] r26_smp_reg,
	output  [47:0] r26_err_reg,
	output  [47:0] r26_idl_reg,
	output  [15:0] r26_lat_reg,
	output  [47:0] r27_smp_reg,
	output  [47:0] r27_err_reg,
	output  [47:0] r27_idl_reg,
	output  [15:0] r27_lat_reg,	
	output  [47:0] r30_smp_reg,
	output  [47:0] r30_err_reg,
	output  [47:0] r30_idl_reg,
	output  [15:0] r30_lat_reg,
	output  [47:0] r31_smp_reg,
	output  [47:0] r31_err_reg,
	output  [47:0] r31_idl_reg,
	output  [15:0] r31_lat_reg,	
	output  [47:0] r32_smp_reg,
	output  [47:0] r32_err_reg,
	output  [47:0] r32_idl_reg,
	output  [15:0] r32_lat_reg,
	output  [47:0] r33_smp_reg,
	output  [47:0] r33_err_reg,
	output  [47:0] r33_idl_reg,
	output  [15:0] r33_lat_reg,
	output  [47:0] r34_smp_reg,
	output  [47:0] r34_err_reg,
	output  [47:0] r34_idl_reg,
	output  [15:0] r34_lat_reg,
	output  [47:0] r35_smp_reg,
	output  [47:0] r35_err_reg,
	output  [47:0] r35_idl_reg,
	output  [15:0] r35_lat_reg,	
	output  [47:0] r36_smp_reg,
	output  [47:0] r36_err_reg,
	output  [47:0] r36_idl_reg,
	output  [15:0] r36_lat_reg,
	output  [47:0] r37_smp_reg,
	output  [47:0] r37_err_reg,
	output  [47:0] r37_idl_reg,
	output  [15:0] r37_lat_reg,
	output  [47:0] r40_smp_reg,
	output  [47:0] r40_err_reg,
	output  [47:0] r40_idl_reg,
	output  [15:0] r40_lat_reg,
	output  [47:0] r41_smp_reg,
	output  [47:0] r41_err_reg,
	output  [47:0] r41_idl_reg,
	output  [15:0] r41_lat_reg,	
	output  [47:0] r42_smp_reg,
	output  [47:0] r42_err_reg,
	output  [47:0] r42_idl_reg,
	output  [15:0] r42_lat_reg,
	output  [47:0] r43_smp_reg,
	output  [47:0] r43_err_reg,
	output  [47:0] r43_idl_reg,
	output  [15:0] r43_lat_reg,
	output  [47:0] r44_smp_reg,
	output  [47:0] r44_err_reg,
	output  [47:0] r44_idl_reg,
	output  [15:0] r44_lat_reg,
	output  [47:0] r45_smp_reg,
	output  [47:0] r45_err_reg,
	output  [47:0] r45_idl_reg,
	output  [15:0] r45_lat_reg,	
	output  [47:0] r46_smp_reg,
	output  [47:0] r46_err_reg,
	output  [47:0] r46_idl_reg,
	output  [15:0] r46_lat_reg,
	output  [47:0] r47_smp_reg,
	output  [47:0] r47_err_reg,
	output  [47:0] r47_idl_reg,
	output  [15:0] r47_lat_reg,
	output  [47:0] r50_smp_reg,
	output  [47:0] r50_err_reg,
	output  [47:0] r50_idl_reg,
	output  [15:0] r50_lat_reg,
	output  [47:0] r51_smp_reg,
	output  [47:0] r51_err_reg,
	output  [47:0] r51_idl_reg,
	output  [15:0] r51_lat_reg,	
	output  [47:0] r52_smp_reg,
	output  [47:0] r52_err_reg,
	output  [47:0] r52_idl_reg,
	output  [15:0] r52_lat_reg,
	output  [47:0] r53_smp_reg,
	output  [47:0] r53_err_reg,
	output  [47:0] r53_idl_reg,
	output  [15:0] r53_lat_reg,
	output  [47:0] r54_smp_reg,
	output  [47:0] r54_err_reg,
	output  [47:0] r54_idl_reg,
	output  [15:0] r54_lat_reg,
	output  [47:0] r55_smp_reg,
	output  [47:0] r55_err_reg,
	output  [47:0] r55_idl_reg,
	output  [15:0] r55_lat_reg,	
	output  [47:0] r56_smp_reg,
	output  [47:0] r56_err_reg,
	output  [47:0] r56_idl_reg,
	output  [15:0] r56_lat_reg,
	output  [47:0] r57_smp_reg,
	output  [47:0] r57_err_reg,
	output  [47:0] r57_idl_reg,
	output  [15:0] r57_lat_reg,	
	output  [47:0] r60_smp_reg,
	output  [47:0] r60_err_reg,
	output  [47:0] r60_idl_reg,
	output  [15:0] r60_lat_reg,
	output  [47:0] r61_smp_reg,
	output  [47:0] r61_err_reg,
	output  [47:0] r61_idl_reg,
	output  [15:0] r61_lat_reg,	
	output  [47:0] r62_smp_reg,
	output  [47:0] r62_err_reg,
	output  [47:0] r62_idl_reg,
	output  [15:0] r62_lat_reg,
	output  [47:0] r63_smp_reg,
	output  [47:0] r63_err_reg,
	output  [47:0] r63_idl_reg,
	output  [15:0] r63_lat_reg,
	output  [47:0] r64_smp_reg,
	output  [47:0] r64_err_reg,
	output  [47:0] r64_idl_reg,
	output  [15:0] r64_lat_reg,
	output  [47:0] r65_smp_reg,
	output  [47:0] r65_err_reg,
	output  [47:0] r65_idl_reg,
	output  [15:0] r65_lat_reg,	
	output  [47:0] r66_smp_reg,
	output  [47:0] r66_err_reg,
	output  [47:0] r66_idl_reg,
	output  [15:0] r66_lat_reg,
	output  [47:0] r67_smp_reg,
	output  [47:0] r67_err_reg,
	output  [47:0] r67_idl_reg,
	output  [15:0] r67_lat_reg,	
	output  [47:0] r70_smp_reg,
	output  [47:0] r70_err_reg,
	output  [47:0] r70_idl_reg,
	output  [15:0] r70_lat_reg,
	output  [47:0] r71_smp_reg,
	output  [47:0] r71_err_reg,
	output  [47:0] r71_idl_reg,
	output  [15:0] r71_lat_reg,	
	output  [47:0] r72_smp_reg,
	output  [47:0] r72_err_reg,
	output  [47:0] r72_idl_reg,
	output  [15:0] r72_lat_reg,
	output  [47:0] r73_smp_reg,
	output  [47:0] r73_err_reg,
	output  [47:0] r73_idl_reg,
	output  [15:0] r73_lat_reg,
	output  [47:0] r74_smp_reg,
	output  [47:0] r74_err_reg,
	output  [47:0] r74_idl_reg,
	output  [15:0] r74_lat_reg,
	output  [47:0] r75_smp_reg,
	output  [47:0] r75_err_reg,
	output  [47:0] r75_idl_reg,
	output  [15:0] r75_lat_reg,	
	output  [47:0] r76_smp_reg,
	output  [47:0] r76_err_reg,
	output  [47:0] r76_idl_reg,
	output  [15:0] r76_lat_reg,
	output  [47:0] r77_smp_reg,
	output  [47:0] r77_err_reg,
	output  [47:0] r77_idl_reg,
	output  [15:0] r77_lat_reg,		
	output  reg   done_stat_reg,
	//----------------------------------
	// aie clock domain
	//----------------------------------	
	input   clk_aie,
	output  test_en_aie,
	input        r00_vld_aie, 
	input [6:0]  r00_smp_aie,
	input [6:0]  r00_err_aie, 
	input [11:0] r00_idl_aie, 
	input [15:0] r00_lat_aie,
	input        r01_vld_aie, 
	input [6:0]  r01_smp_aie,
	input [6:0]  r01_err_aie, 
	input [11:0] r01_idl_aie, 
	input [15:0] r01_lat_aie,
	input        r02_vld_aie, 
	input [6:0]  r02_smp_aie,
	input [6:0]  r02_err_aie, 
	input [11:0] r02_idl_aie, 
	input [15:0] r02_lat_aie,
	input        r03_vld_aie, 
	input [6:0]  r03_smp_aie,
	input [6:0]  r03_err_aie, 
	input [11:0] r03_idl_aie, 
	input [15:0] r03_lat_aie,
	input        r04_vld_aie, 
	input [6:0]  r04_smp_aie,
	input [6:0]  r04_err_aie, 
	input [11:0] r04_idl_aie, 
	input [15:0] r04_lat_aie,
	input        r05_vld_aie, 
	input [6:0]  r05_smp_aie,
	input [6:0]  r05_err_aie, 
	input [11:0] r05_idl_aie, 
	input [15:0] r05_lat_aie,
	input        r06_vld_aie, 
	input [6:0]  r06_smp_aie,
	input [6:0]  r06_err_aie, 
	input [11:0] r06_idl_aie, 
	input [15:0] r06_lat_aie,
	input        r07_vld_aie, 
	input [6:0]  r07_smp_aie,
	input [6:0]  r07_err_aie, 
	input [11:0] r07_idl_aie, 
	input [15:0] r07_lat_aie,
	input        r10_vld_aie, 
	input [6:0]  r10_smp_aie,
	input [6:0]  r10_err_aie, 
	input [11:0] r10_idl_aie, 
	input [15:0] r10_lat_aie,
	input        r11_vld_aie, 
	input [6:0]  r11_smp_aie,
	input [6:0]  r11_err_aie, 
	input [11:0] r11_idl_aie, 
	input [15:0] r11_lat_aie,
	input        r12_vld_aie, 
	input [6:0]  r12_smp_aie,
	input [6:0]  r12_err_aie, 
	input [11:0] r12_idl_aie, 
	input [15:0] r12_lat_aie,
	input        r13_vld_aie, 
	input [6:0]  r13_smp_aie,
	input [6:0]  r13_err_aie, 
	input [11:0] r13_idl_aie, 
	input [15:0] r13_lat_aie,
	input        r14_vld_aie, 
	input [6:0]  r14_smp_aie,
	input [6:0]  r14_err_aie, 
	input [11:0] r14_idl_aie, 
	input [15:0] r14_lat_aie,
	input        r15_vld_aie, 
	input [6:0]  r15_smp_aie,
	input [6:0]  r15_err_aie, 
	input [11:0] r15_idl_aie, 
	input [15:0] r15_lat_aie,
	input        r16_vld_aie, 
	input [6:0]  r16_smp_aie,
	input [6:0]  r16_err_aie, 
	input [11:0] r16_idl_aie, 
	input [15:0] r16_lat_aie,
	input        r17_vld_aie, 
	input [6:0]  r17_smp_aie,
	input [6:0]  r17_err_aie, 
	input [11:0] r17_idl_aie, 
	input [15:0] r17_lat_aie,
	input        r20_vld_aie, 
	input [6:0]  r20_smp_aie,
	input [6:0]  r20_err_aie, 
	input [11:0] r20_idl_aie, 
	input [15:0] r20_lat_aie,
	input        r21_vld_aie, 
	input [6:0]  r21_smp_aie,
	input [6:0]  r21_err_aie, 
	input [11:0] r21_idl_aie, 
	input [15:0] r21_lat_aie,
	input        r22_vld_aie, 
	input [6:0]  r22_smp_aie,
	input [6:0]  r22_err_aie, 
	input [11:0] r22_idl_aie, 
	input [15:0] r22_lat_aie,
	input        r23_vld_aie, 
	input [6:0]  r23_smp_aie,
	input [6:0]  r23_err_aie, 
	input [11:0] r23_idl_aie, 
	input [15:0] r23_lat_aie,
	input        r24_vld_aie, 
	input [6:0]  r24_smp_aie,
	input [6:0]  r24_err_aie, 
	input [11:0] r24_idl_aie, 
	input [15:0] r24_lat_aie,
	input        r25_vld_aie, 
	input [6:0]  r25_smp_aie,
	input [6:0]  r25_err_aie, 
	input [11:0] r25_idl_aie, 
	input [15:0] r25_lat_aie,
	input        r26_vld_aie, 
	input [6:0]  r26_smp_aie,
	input [6:0]  r26_err_aie, 
	input [11:0] r26_idl_aie, 
	input [15:0] r26_lat_aie,
	input        r27_vld_aie, 
	input [6:0]  r27_smp_aie,
	input [6:0]  r27_err_aie, 
	input [11:0] r27_idl_aie, 
	input [15:0] r27_lat_aie,
	input        r30_vld_aie, 
	input [6:0]  r30_smp_aie,
	input [6:0]  r30_err_aie, 
	input [11:0] r30_idl_aie, 
	input [15:0] r30_lat_aie,
	input        r31_vld_aie, 
	input [6:0]  r31_smp_aie,
	input [6:0]  r31_err_aie, 
	input [11:0] r31_idl_aie, 
	input [15:0] r31_lat_aie,
	input        r32_vld_aie, 
	input [6:0]  r32_smp_aie,
	input [6:0]  r32_err_aie, 
	input [11:0] r32_idl_aie, 
	input [15:0] r32_lat_aie,
	input        r33_vld_aie, 
	input [6:0]  r33_smp_aie,
	input [6:0]  r33_err_aie, 
	input [11:0] r33_idl_aie, 
	input [15:0] r33_lat_aie,
	input        r34_vld_aie, 
	input [6:0]  r34_smp_aie,
	input [6:0]  r34_err_aie, 
	input [11:0] r34_idl_aie, 
	input [15:0] r34_lat_aie,
	input        r35_vld_aie, 
	input [6:0]  r35_smp_aie,
	input [6:0]  r35_err_aie, 
	input [11:0] r35_idl_aie, 
	input [15:0] r35_lat_aie,
	input        r36_vld_aie, 
	input [6:0]  r36_smp_aie,
	input [6:0]  r36_err_aie, 
	input [11:0] r36_idl_aie, 
	input [15:0] r36_lat_aie,
	input        r37_vld_aie, 
	input [6:0]  r37_smp_aie,
	input [6:0]  r37_err_aie, 
	input [11:0] r37_idl_aie, 
	input [15:0] r37_lat_aie,
	input        r40_vld_aie, 
	input [6:0]  r40_smp_aie,
	input [6:0]  r40_err_aie, 
	input [11:0] r40_idl_aie, 
	input [15:0] r40_lat_aie,
	input        r41_vld_aie, 
	input [6:0]  r41_smp_aie,
	input [6:0]  r41_err_aie, 
	input [11:0] r41_idl_aie, 
	input [15:0] r41_lat_aie,
	input        r42_vld_aie, 
	input [6:0]  r42_smp_aie,
	input [6:0]  r42_err_aie, 
	input [11:0] r42_idl_aie, 
	input [15:0] r42_lat_aie,
	input        r43_vld_aie, 
	input [6:0]  r43_smp_aie,
	input [6:0]  r43_err_aie, 
	input [11:0] r43_idl_aie, 
	input [15:0] r43_lat_aie,
	input        r44_vld_aie, 
	input [6:0]  r44_smp_aie,
	input [6:0]  r44_err_aie, 
	input [11:0] r44_idl_aie, 
	input [15:0] r44_lat_aie,
	input        r45_vld_aie, 
	input [6:0]  r45_smp_aie,
	input [6:0]  r45_err_aie, 
	input [11:0] r45_idl_aie, 
	input [15:0] r45_lat_aie,
	input        r46_vld_aie, 
	input [6:0]  r46_smp_aie,
	input [6:0]  r46_err_aie, 
	input [11:0] r46_idl_aie, 
	input [15:0] r46_lat_aie,
	input        r47_vld_aie, 
	input [6:0]  r47_smp_aie,
	input [6:0]  r47_err_aie, 
	input [11:0] r47_idl_aie, 
	input [15:0] r47_lat_aie,
	input        r50_vld_aie, 
	input [6:0]  r50_smp_aie,
	input [6:0]  r50_err_aie, 
	input [11:0] r50_idl_aie, 
	input [15:0] r50_lat_aie,
	input        r51_vld_aie, 
	input [6:0]  r51_smp_aie,
	input [6:0]  r51_err_aie, 
	input [11:0] r51_idl_aie, 
	input [15:0] r51_lat_aie,
	input        r52_vld_aie, 
	input [6:0]  r52_smp_aie,
	input [6:0]  r52_err_aie, 
	input [11:0] r52_idl_aie, 
	input [15:0] r52_lat_aie,
	input        r53_vld_aie, 
	input [6:0]  r53_smp_aie,
	input [6:0]  r53_err_aie, 
	input [11:0] r53_idl_aie, 
	input [15:0] r53_lat_aie,
	input        r54_vld_aie, 
	input [6:0]  r54_smp_aie,
	input [6:0]  r54_err_aie, 
	input [11:0] r54_idl_aie, 
	input [15:0] r54_lat_aie,
	input        r55_vld_aie, 
	input [6:0]  r55_smp_aie,
	input [6:0]  r55_err_aie, 
	input [11:0] r55_idl_aie, 
	input [15:0] r55_lat_aie,
	input        r56_vld_aie, 
	input [6:0]  r56_smp_aie,
	input [6:0]  r56_err_aie, 
	input [11:0] r56_idl_aie, 
	input [15:0] r56_lat_aie,
	input        r57_vld_aie, 
	input [6:0]  r57_smp_aie,
	input [6:0]  r57_err_aie, 
	input [11:0] r57_idl_aie, 
	input [15:0] r57_lat_aie,
	input        r60_vld_aie, 
	input [6:0]  r60_smp_aie,
	input [6:0]  r60_err_aie, 
	input [11:0] r60_idl_aie, 
	input [15:0] r60_lat_aie,
	input        r61_vld_aie, 
	input [6:0]  r61_smp_aie,
	input [6:0]  r61_err_aie, 
	input [11:0] r61_idl_aie, 
	input [15:0] r61_lat_aie,
	input        r62_vld_aie, 
	input [6:0]  r62_smp_aie,
	input [6:0]  r62_err_aie, 
	input [11:0] r62_idl_aie, 
	input [15:0] r62_lat_aie,
	input        r63_vld_aie, 
	input [6:0]  r63_smp_aie,
	input [6:0]  r63_err_aie, 
	input [11:0] r63_idl_aie, 
	input [15:0] r63_lat_aie,
	input        r64_vld_aie, 
	input [6:0]  r64_smp_aie,
	input [6:0]  r64_err_aie, 
	input [11:0] r64_idl_aie, 
	input [15:0] r64_lat_aie,
	input        r65_vld_aie, 
	input [6:0]  r65_smp_aie,
	input [6:0]  r65_err_aie, 
	input [11:0] r65_idl_aie, 
	input [15:0] r65_lat_aie,
	input        r66_vld_aie, 
	input [6:0]  r66_smp_aie,
	input [6:0]  r66_err_aie, 
	input [11:0] r66_idl_aie, 
	input [15:0] r66_lat_aie,
	input        r67_vld_aie, 
	input [6:0]  r67_smp_aie,
	input [6:0]  r67_err_aie, 
	input [11:0] r67_idl_aie, 
	input [15:0] r67_lat_aie,
	input        r70_vld_aie, 
	input [6:0]  r70_smp_aie,
	input [6:0]  r70_err_aie, 
	input [11:0] r70_idl_aie, 
	input [15:0] r70_lat_aie,
	input        r71_vld_aie, 
	input [6:0]  r71_smp_aie,
	input [6:0]  r71_err_aie, 
	input [11:0] r71_idl_aie, 
	input [15:0] r71_lat_aie,
	input        r72_vld_aie, 
	input [6:0]  r72_smp_aie,
	input [6:0]  r72_err_aie, 
	input [11:0] r72_idl_aie, 
	input [15:0] r72_lat_aie,
	input        r73_vld_aie, 
	input [6:0]  r73_smp_aie,
	input [6:0]  r73_err_aie, 
	input [11:0] r73_idl_aie, 
	input [15:0] r73_lat_aie,
	input        r74_vld_aie, 
	input [6:0]  r74_smp_aie,
	input [6:0]  r74_err_aie, 
	input [11:0] r74_idl_aie, 
	input [15:0] r74_lat_aie,
	input        r75_vld_aie, 
	input [6:0]  r75_smp_aie,
	input [6:0]  r75_err_aie, 
	input [11:0] r75_idl_aie, 
	input [15:0] r75_lat_aie,
	input        r76_vld_aie, 
	input [6:0]  r76_smp_aie,
	input [6:0]  r76_err_aie, 
	input [11:0] r76_idl_aie, 
	input [15:0] r76_lat_aie,
	input        r77_vld_aie, 
	input [6:0]  r77_smp_aie,
	input [6:0]  r77_err_aie, 
	input [11:0] r77_idl_aie, 
	input [15:0] r77_lat_aie,		
	input [63:0] done_aie
);

wire [63:0] s_done;
reg test_en_s;

//----------------------------------------
// REG -> AIE
//----------------------------------------
xpm_cdc_single #(
 .DEST_SYNC_FF(4), // DECIMAL; range: 2-10
 .INIT_SYNC_FF(1), // DECIMAL; 0=disable simulation init values, 1=enable simulation init values
 .SIM_ASSERT_CHK(0), // DECIMAL; 0=disable simulation messages, 1=enable simulation messages
 .SRC_INPUT_REG(0) // DECIMAL; 0=do not register input, 1=register input
)
CDC0(
 .dest_out(test_en_aie), // 1-bit output: src_in synchronized to the destination clock domain. This output is
 // registered.
 .dest_clk(clk_aie), // 1-bit input: Clock signal for the destination clock domain.
 .src_clk(), // 1-bit input: optional; required when SRC_INPUT_REG = 1
 .src_in(test_en_reg) // 1-bit input: Input signal to be synchronized to dest_clk domain.
);


always @(posedge clk_reg) done_stat_reg <= &s_done;
always @(posedge clk_reg) test_en_s <= test_en_reg;

//----------------------------------------
// Test Result Registers
//----------------------------------------
tst_dout_xclk_results R00(clk_reg, test_en_s, r00_vld_aie, r00_smp_aie, r00_err_aie, r00_idl_aie, r00_lat_aie, done_aie[ 0],	r00_smp_reg, r00_err_reg, r00_idl_reg, r00_lat_reg, s_done[ 0]);
tst_dout_xclk_results R01(clk_reg, test_en_s, r01_vld_aie, r01_smp_aie, r01_err_aie, r01_idl_aie, r01_lat_aie, done_aie[ 1],	r01_smp_reg, r01_err_reg, r01_idl_reg, r01_lat_reg, s_done[ 1]);
tst_dout_xclk_results R02(clk_reg, test_en_s, r02_vld_aie, r02_smp_aie, r02_err_aie, r02_idl_aie, r02_lat_aie, done_aie[ 2],	r02_smp_reg, r02_err_reg, r02_idl_reg, r02_lat_reg, s_done[ 2]);
tst_dout_xclk_results R03(clk_reg, test_en_s, r03_vld_aie, r03_smp_aie, r03_err_aie, r03_idl_aie, r03_lat_aie, done_aie[ 3],	r03_smp_reg, r03_err_reg, r03_idl_reg, r03_lat_reg, s_done[ 3]);
tst_dout_xclk_results R04(clk_reg, test_en_s, r04_vld_aie, r04_smp_aie, r04_err_aie, r04_idl_aie, r04_lat_aie, done_aie[ 4],	r04_smp_reg, r04_err_reg, r04_idl_reg, r04_lat_reg, s_done[ 4]);
tst_dout_xclk_results R05(clk_reg, test_en_s, r05_vld_aie, r05_smp_aie, r05_err_aie, r05_idl_aie, r05_lat_aie, done_aie[ 5],	r05_smp_reg, r05_err_reg, r05_idl_reg, r05_lat_reg, s_done[ 5]);
tst_dout_xclk_results R06(clk_reg, test_en_s, r06_vld_aie, r06_smp_aie, r06_err_aie, r06_idl_aie, r06_lat_aie, done_aie[ 6],	r06_smp_reg, r06_err_reg, r06_idl_reg, r06_lat_reg, s_done[ 6]);
tst_dout_xclk_results R07(clk_reg, test_en_s, r07_vld_aie, r07_smp_aie, r07_err_aie, r07_idl_aie, r07_lat_aie, done_aie[ 7],	r07_smp_reg, r07_err_reg, r07_idl_reg, r07_lat_reg, s_done[ 7]);
tst_dout_xclk_results R10(clk_reg, test_en_s, r10_vld_aie, r10_smp_aie, r10_err_aie, r10_idl_aie, r10_lat_aie, done_aie[8+0],	r10_smp_reg, r10_err_reg, r10_idl_reg, r10_lat_reg, s_done[8+0]);
tst_dout_xclk_results R11(clk_reg, test_en_s, r11_vld_aie, r11_smp_aie, r11_err_aie, r11_idl_aie, r11_lat_aie, done_aie[8+1],	r11_smp_reg, r11_err_reg, r11_idl_reg, r11_lat_reg, s_done[8+1]);
tst_dout_xclk_results R12(clk_reg, test_en_s, r12_vld_aie, r12_smp_aie, r12_err_aie, r12_idl_aie, r12_lat_aie, done_aie[8+2],	r12_smp_reg, r12_err_reg, r12_idl_reg, r12_lat_reg, s_done[8+2]);
tst_dout_xclk_results R13(clk_reg, test_en_s, r13_vld_aie, r13_smp_aie, r13_err_aie, r13_idl_aie, r13_lat_aie, done_aie[8+3],	r13_smp_reg, r13_err_reg, r13_idl_reg, r13_lat_reg, s_done[8+3]);
tst_dout_xclk_results R14(clk_reg, test_en_s, r14_vld_aie, r14_smp_aie, r14_err_aie, r14_idl_aie, r14_lat_aie, done_aie[8+4],	r14_smp_reg, r14_err_reg, r14_idl_reg, r14_lat_reg, s_done[8+4]);
tst_dout_xclk_results R15(clk_reg, test_en_s, r15_vld_aie, r15_smp_aie, r15_err_aie, r15_idl_aie, r15_lat_aie, done_aie[8+5],	r15_smp_reg, r15_err_reg, r15_idl_reg, r15_lat_reg, s_done[8+5]);
tst_dout_xclk_results R16(clk_reg, test_en_s, r16_vld_aie, r16_smp_aie, r16_err_aie, r16_idl_aie, r16_lat_aie, done_aie[8+6],	r16_smp_reg, r16_err_reg, r16_idl_reg, r16_lat_reg, s_done[8+6]);
tst_dout_xclk_results R17(clk_reg, test_en_s, r17_vld_aie, r17_smp_aie, r17_err_aie, r17_idl_aie, r17_lat_aie, done_aie[8+7],	r17_smp_reg, r17_err_reg, r17_idl_reg, r17_lat_reg, s_done[8+7]);
tst_dout_xclk_results R20(clk_reg, test_en_s, r20_vld_aie, r20_smp_aie, r20_err_aie, r20_idl_aie, r20_lat_aie, done_aie[8*2+0],	r20_smp_reg, r20_err_reg, r20_idl_reg, r20_lat_reg, s_done[8*2+0]);
tst_dout_xclk_results R21(clk_reg, test_en_s, r21_vld_aie, r21_smp_aie, r21_err_aie, r21_idl_aie, r21_lat_aie, done_aie[8*2+1],	r21_smp_reg, r21_err_reg, r21_idl_reg, r21_lat_reg, s_done[8*2+1]);
tst_dout_xclk_results R22(clk_reg, test_en_s, r22_vld_aie, r22_smp_aie, r22_err_aie, r22_idl_aie, r22_lat_aie, done_aie[8*2+2],	r22_smp_reg, r22_err_reg, r22_idl_reg, r22_lat_reg, s_done[8*2+2]);
tst_dout_xclk_results R23(clk_reg, test_en_s, r23_vld_aie, r23_smp_aie, r23_err_aie, r23_idl_aie, r23_lat_aie, done_aie[8*2+3],	r23_smp_reg, r23_err_reg, r23_idl_reg, r23_lat_reg, s_done[8*2+3]);
tst_dout_xclk_results R24(clk_reg, test_en_s, r24_vld_aie, r24_smp_aie, r24_err_aie, r24_idl_aie, r24_lat_aie, done_aie[8*2+4],	r24_smp_reg, r24_err_reg, r24_idl_reg, r24_lat_reg, s_done[8*2+4]);
tst_dout_xclk_results R25(clk_reg, test_en_s, r25_vld_aie, r25_smp_aie, r25_err_aie, r25_idl_aie, r25_lat_aie, done_aie[8*2+5],	r25_smp_reg, r25_err_reg, r25_idl_reg, r25_lat_reg, s_done[8*2+5]);
tst_dout_xclk_results R26(clk_reg, test_en_s, r26_vld_aie, r26_smp_aie, r26_err_aie, r26_idl_aie, r26_lat_aie, done_aie[8*2+6],	r26_smp_reg, r26_err_reg, r26_idl_reg, r26_lat_reg, s_done[8*2+6]);
tst_dout_xclk_results R27(clk_reg, test_en_s, r27_vld_aie, r27_smp_aie, r27_err_aie, r27_idl_aie, r27_lat_aie, done_aie[8*2+7],	r27_smp_reg, r27_err_reg, r27_idl_reg, r27_lat_reg, s_done[8*2+7]);
tst_dout_xclk_results R30(clk_reg, test_en_s, r30_vld_aie, r30_smp_aie, r30_err_aie, r30_idl_aie, r30_lat_aie, done_aie[8*3+0],	r30_smp_reg, r30_err_reg, r30_idl_reg, r30_lat_reg, s_done[8*3+0]);
tst_dout_xclk_results R31(clk_reg, test_en_s, r31_vld_aie, r31_smp_aie, r31_err_aie, r31_idl_aie, r31_lat_aie, done_aie[8*3+1],	r31_smp_reg, r31_err_reg, r31_idl_reg, r31_lat_reg, s_done[8*3+1]);
tst_dout_xclk_results R32(clk_reg, test_en_s, r32_vld_aie, r32_smp_aie, r32_err_aie, r32_idl_aie, r32_lat_aie, done_aie[8*3+2],	r32_smp_reg, r32_err_reg, r32_idl_reg, r32_lat_reg, s_done[8*3+2]);
tst_dout_xclk_results R33(clk_reg, test_en_s, r33_vld_aie, r33_smp_aie, r33_err_aie, r33_idl_aie, r33_lat_aie, done_aie[8*3+3],	r33_smp_reg, r33_err_reg, r33_idl_reg, r33_lat_reg, s_done[8*3+3]);
tst_dout_xclk_results R34(clk_reg, test_en_s, r34_vld_aie, r34_smp_aie, r34_err_aie, r34_idl_aie, r34_lat_aie, done_aie[8*3+4],	r34_smp_reg, r34_err_reg, r34_idl_reg, r34_lat_reg, s_done[8*3+4]);
tst_dout_xclk_results R35(clk_reg, test_en_s, r35_vld_aie, r35_smp_aie, r35_err_aie, r35_idl_aie, r35_lat_aie, done_aie[8*3+5],	r35_smp_reg, r35_err_reg, r35_idl_reg, r35_lat_reg, s_done[8*3+5]);
tst_dout_xclk_results R36(clk_reg, test_en_s, r36_vld_aie, r36_smp_aie, r36_err_aie, r36_idl_aie, r36_lat_aie, done_aie[8*3+6],	r36_smp_reg, r36_err_reg, r36_idl_reg, r36_lat_reg, s_done[8*3+6]);
tst_dout_xclk_results R37(clk_reg, test_en_s, r37_vld_aie, r37_smp_aie, r37_err_aie, r37_idl_aie, r37_lat_aie, done_aie[8*3+7],	r37_smp_reg, r37_err_reg, r37_idl_reg, r37_lat_reg, s_done[8*3+7]);
tst_dout_xclk_results R40(clk_reg, test_en_s, r40_vld_aie, r40_smp_aie, r40_err_aie, r40_idl_aie, r40_lat_aie, done_aie[8*4+0],	r40_smp_reg, r40_err_reg, r40_idl_reg, r40_lat_reg, s_done[8*4+0]);
tst_dout_xclk_results R41(clk_reg, test_en_s, r41_vld_aie, r41_smp_aie, r41_err_aie, r41_idl_aie, r41_lat_aie, done_aie[8*4+1],	r41_smp_reg, r41_err_reg, r41_idl_reg, r41_lat_reg, s_done[8*4+1]);
tst_dout_xclk_results R42(clk_reg, test_en_s, r42_vld_aie, r42_smp_aie, r42_err_aie, r42_idl_aie, r42_lat_aie, done_aie[8*4+2],	r42_smp_reg, r42_err_reg, r42_idl_reg, r42_lat_reg, s_done[8*4+2]);
tst_dout_xclk_results R43(clk_reg, test_en_s, r43_vld_aie, r43_smp_aie, r43_err_aie, r43_idl_aie, r43_lat_aie, done_aie[8*4+3],	r43_smp_reg, r43_err_reg, r43_idl_reg, r43_lat_reg, s_done[8*4+3]);
tst_dout_xclk_results R44(clk_reg, test_en_s, r44_vld_aie, r44_smp_aie, r44_err_aie, r44_idl_aie, r44_lat_aie, done_aie[8*4+4],	r44_smp_reg, r44_err_reg, r44_idl_reg, r44_lat_reg, s_done[8*4+4]);
tst_dout_xclk_results R45(clk_reg, test_en_s, r45_vld_aie, r45_smp_aie, r45_err_aie, r45_idl_aie, r45_lat_aie, done_aie[8*4+5],	r45_smp_reg, r45_err_reg, r45_idl_reg, r45_lat_reg, s_done[8*4+5]);
tst_dout_xclk_results R46(clk_reg, test_en_s, r46_vld_aie, r46_smp_aie, r46_err_aie, r46_idl_aie, r46_lat_aie, done_aie[8*4+6],	r46_smp_reg, r46_err_reg, r46_idl_reg, r46_lat_reg, s_done[8*4+6]);
tst_dout_xclk_results R47(clk_reg, test_en_s, r47_vld_aie, r47_smp_aie, r47_err_aie, r47_idl_aie, r47_lat_aie, done_aie[8*4+7],	r47_smp_reg, r47_err_reg, r47_idl_reg, r47_lat_reg, s_done[8*4+7]);
tst_dout_xclk_results R50(clk_reg, test_en_s, r50_vld_aie, r50_smp_aie, r50_err_aie, r50_idl_aie, r50_lat_aie, done_aie[8*5+0],	r50_smp_reg, r50_err_reg, r50_idl_reg, r50_lat_reg, s_done[8*5+0]);
tst_dout_xclk_results R51(clk_reg, test_en_s, r51_vld_aie, r51_smp_aie, r51_err_aie, r51_idl_aie, r51_lat_aie, done_aie[8*5+1],	r51_smp_reg, r51_err_reg, r51_idl_reg, r51_lat_reg, s_done[8*5+1]);
tst_dout_xclk_results R52(clk_reg, test_en_s, r52_vld_aie, r52_smp_aie, r52_err_aie, r52_idl_aie, r52_lat_aie, done_aie[8*5+2],	r52_smp_reg, r52_err_reg, r52_idl_reg, r52_lat_reg, s_done[8*5+2]);
tst_dout_xclk_results R53(clk_reg, test_en_s, r53_vld_aie, r53_smp_aie, r53_err_aie, r53_idl_aie, r53_lat_aie, done_aie[8*5+3],	r53_smp_reg, r53_err_reg, r53_idl_reg, r53_lat_reg, s_done[8*5+3]);
tst_dout_xclk_results R54(clk_reg, test_en_s, r54_vld_aie, r54_smp_aie, r54_err_aie, r54_idl_aie, r54_lat_aie, done_aie[8*5+4],	r54_smp_reg, r54_err_reg, r54_idl_reg, r54_lat_reg, s_done[8*5+4]);
tst_dout_xclk_results R55(clk_reg, test_en_s, r55_vld_aie, r55_smp_aie, r55_err_aie, r55_idl_aie, r55_lat_aie, done_aie[8*5+5],	r55_smp_reg, r55_err_reg, r55_idl_reg, r55_lat_reg, s_done[8*5+5]);
tst_dout_xclk_results R56(clk_reg, test_en_s, r56_vld_aie, r56_smp_aie, r56_err_aie, r56_idl_aie, r56_lat_aie, done_aie[8*5+6],	r56_smp_reg, r56_err_reg, r56_idl_reg, r56_lat_reg, s_done[8*5+6]);
tst_dout_xclk_results R57(clk_reg, test_en_s, r57_vld_aie, r57_smp_aie, r57_err_aie, r57_idl_aie, r57_lat_aie, done_aie[8*5+7],	r57_smp_reg, r57_err_reg, r57_idl_reg, r57_lat_reg, s_done[8*5+7]);
tst_dout_xclk_results R60(clk_reg, test_en_s, r60_vld_aie, r60_smp_aie, r60_err_aie, r60_idl_aie, r60_lat_aie, done_aie[8*6+0],	r60_smp_reg, r60_err_reg, r60_idl_reg, r60_lat_reg, s_done[8*6+0]);
tst_dout_xclk_results R61(clk_reg, test_en_s, r61_vld_aie, r61_smp_aie, r61_err_aie, r61_idl_aie, r61_lat_aie, done_aie[8*6+1],	r61_smp_reg, r61_err_reg, r61_idl_reg, r61_lat_reg, s_done[8*6+1]);
tst_dout_xclk_results R62(clk_reg, test_en_s, r62_vld_aie, r62_smp_aie, r62_err_aie, r62_idl_aie, r62_lat_aie, done_aie[8*6+2],	r62_smp_reg, r62_err_reg, r62_idl_reg, r62_lat_reg, s_done[8*6+2]);
tst_dout_xclk_results R63(clk_reg, test_en_s, r63_vld_aie, r63_smp_aie, r63_err_aie, r63_idl_aie, r63_lat_aie, done_aie[8*6+3],	r63_smp_reg, r63_err_reg, r63_idl_reg, r63_lat_reg, s_done[8*6+3]);
tst_dout_xclk_results R64(clk_reg, test_en_s, r64_vld_aie, r64_smp_aie, r64_err_aie, r64_idl_aie, r64_lat_aie, done_aie[8*6+4],	r64_smp_reg, r64_err_reg, r64_idl_reg, r64_lat_reg, s_done[8*6+4]);
tst_dout_xclk_results R65(clk_reg, test_en_s, r65_vld_aie, r65_smp_aie, r65_err_aie, r65_idl_aie, r65_lat_aie, done_aie[8*6+5],	r65_smp_reg, r65_err_reg, r65_idl_reg, r65_lat_reg, s_done[8*6+5]);
tst_dout_xclk_results R66(clk_reg, test_en_s, r66_vld_aie, r66_smp_aie, r66_err_aie, r66_idl_aie, r66_lat_aie, done_aie[8*6+6],	r66_smp_reg, r66_err_reg, r66_idl_reg, r66_lat_reg, s_done[8*6+6]);
tst_dout_xclk_results R67(clk_reg, test_en_s, r67_vld_aie, r67_smp_aie, r67_err_aie, r67_idl_aie, r67_lat_aie, done_aie[8*6+7],	r67_smp_reg, r67_err_reg, r67_idl_reg, r67_lat_reg, s_done[8*6+7]);
tst_dout_xclk_results R70(clk_reg, test_en_s, r70_vld_aie, r70_smp_aie, r70_err_aie, r70_idl_aie, r70_lat_aie, done_aie[8*7+0],	r70_smp_reg, r70_err_reg, r70_idl_reg, r70_lat_reg, s_done[8*7+0]);
tst_dout_xclk_results R71(clk_reg, test_en_s, r71_vld_aie, r71_smp_aie, r71_err_aie, r71_idl_aie, r71_lat_aie, done_aie[8*7+1],	r71_smp_reg, r71_err_reg, r71_idl_reg, r71_lat_reg, s_done[8*7+1]);
tst_dout_xclk_results R72(clk_reg, test_en_s, r72_vld_aie, r72_smp_aie, r72_err_aie, r72_idl_aie, r72_lat_aie, done_aie[8*7+2],	r72_smp_reg, r72_err_reg, r72_idl_reg, r72_lat_reg, s_done[8*7+2]);
tst_dout_xclk_results R73(clk_reg, test_en_s, r73_vld_aie, r73_smp_aie, r73_err_aie, r73_idl_aie, r73_lat_aie, done_aie[8*7+3],	r73_smp_reg, r73_err_reg, r73_idl_reg, r73_lat_reg, s_done[8*7+3]);
tst_dout_xclk_results R74(clk_reg, test_en_s, r74_vld_aie, r74_smp_aie, r74_err_aie, r74_idl_aie, r74_lat_aie, done_aie[8*7+4],	r74_smp_reg, r74_err_reg, r74_idl_reg, r74_lat_reg, s_done[8*7+4]);
tst_dout_xclk_results R75(clk_reg, test_en_s, r75_vld_aie, r75_smp_aie, r75_err_aie, r75_idl_aie, r75_lat_aie, done_aie[8*7+5],	r75_smp_reg, r75_err_reg, r75_idl_reg, r75_lat_reg, s_done[8*7+5]);
tst_dout_xclk_results R76(clk_reg, test_en_s, r76_vld_aie, r76_smp_aie, r76_err_aie, r76_idl_aie, r76_lat_aie, done_aie[8*7+6],	r76_smp_reg, r76_err_reg, r76_idl_reg, r76_lat_reg, s_done[8*7+6]);
tst_dout_xclk_results R77(clk_reg, test_en_s, r77_vld_aie, r77_smp_aie, r77_err_aie, r77_idl_aie, r77_lat_aie, done_aie[8*7+7],	r77_smp_reg, r77_err_reg, r77_idl_reg, r77_lat_reg, s_done[8*7+7]);


endmodule
